
module SECBADAEC_encoder(input [127:0] message, output [135:0] codeword);

	assign codeword[135:8] = message[127:0];
	assign codeword[7] = ^(message&128'b11011001001011010101010111011010010001110010001000100100001010011110101101000010010001011001000101111110100000100101111111001100);
	assign codeword[6] = ^(message&128'b10110011010110101010101110110100100011100100010001001000010100111101011110000101100010110010001111111101000001001011111010011000);
	assign codeword[5] = ^(message&128'b10111110100110000000001010110011010110101010101110110100100011100100010001001000010100111101011110000101100010110010001111111101);
	assign codeword[4] = ^(message&128'b10100101000111000101000010111101111100100111010101001101001101000110001011010010111000100011111001110100100101000001100100110111);
	assign codeword[3] = ^(message&128'b01001011001110011010000001111011111001011110101010011011011010001100010010100100110001010111110111101000001010000011001001101111);
	assign codeword[2] = ^(message&128'b10010111011100110100000011110110110010111101010100110110110100011000100001001001100010101111101011010000010100010110010011011111);
	assign codeword[1] = ^(message&128'b11110110110010111101010100110110110100011000100001001001100010101111101011010000010100010110010011011111001000001001011101110011);
	assign codeword[0] = ^(message&128'b11101100100101101010101001101101101000110001000110010010000101001111010110100001101000101100100010111111010000010010111111100110);

endmodule

